module Input_Device_module(Data_in, Data_out);
    input [31:0]Data_in;
    output [31:0]Data_out;
    
    assign Data_out = Data_in;
endmodule
